// alarm.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module alarm (
		output wire        alarm_export,    //    alarm.export
		input  wire [3:0]  buttons_export,  //  buttons.export
		input  wire        clk_clk,         //      clk.clk
		output wire [15:0] hours_export,    //    hours.export
		output wire [9:0]  leds_export,     //     leds.export
		output wire [15:0] minutes_export,  //  minutes.export
		input  wire        reset_reset_n,   //    reset.reset_n
		output wire [15:0] seconds_export,  //  seconds.export
		input  wire [1:0]  switches_export, // switches.export
		input  wire        uart_RXD,        //     uart.RXD
		output wire        uart_TXD         //         .TXD
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [18:0] cpu_data_master_address;                              // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                 // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [18:0] cpu_instruction_master_address;                       // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                          // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire         mm_interconnect_0_uart_avalon_rs232_slave_chipselect; // mm_interconnect_0:UART_avalon_rs232_slave_chipselect -> UART:chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_rs232_slave_readdata;   // UART:readdata -> mm_interconnect_0:UART_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_uart_avalon_rs232_slave_address;    // mm_interconnect_0:UART_avalon_rs232_slave_address -> UART:address
	wire         mm_interconnect_0_uart_avalon_rs232_slave_read;       // mm_interconnect_0:UART_avalon_rs232_slave_read -> UART:read
	wire   [3:0] mm_interconnect_0_uart_avalon_rs232_slave_byteenable; // mm_interconnect_0:UART_avalon_rs232_slave_byteenable -> UART:byteenable
	wire         mm_interconnect_0_uart_avalon_rs232_slave_write;      // mm_interconnect_0:UART_avalon_rs232_slave_write -> UART:write
	wire  [31:0] mm_interconnect_0_uart_avalon_rs232_slave_writedata;  // mm_interconnect_0:UART_avalon_rs232_slave_writedata -> UART:writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;       // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;        // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [12:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_rom_s1_chipselect;                  // mm_interconnect_0:ROM_s1_chipselect -> ROM:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                    // ROM:readdata -> mm_interconnect_0:ROM_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                 // mm_interconnect_0:ROM_s1_debugaccess -> ROM:debugaccess
	wire  [14:0] mm_interconnect_0_rom_s1_address;                     // mm_interconnect_0:ROM_s1_address -> ROM:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                  // mm_interconnect_0:ROM_s1_byteenable -> ROM:byteenable
	wire         mm_interconnect_0_rom_s1_write;                       // mm_interconnect_0:ROM_s1_write -> ROM:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                   // mm_interconnect_0:ROM_s1_writedata -> ROM:writedata
	wire         mm_interconnect_0_rom_s1_clken;                       // mm_interconnect_0:ROM_s1_clken -> ROM:clken
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                // BUTTONS:readdata -> mm_interconnect_0:BUTTONS_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                 // mm_interconnect_0:BUTTONS_s1_address -> BUTTONS:address
	wire         mm_interconnect_0_leds_s1_chipselect;                 // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                   // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                    // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                      // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                  // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_seconds_s1_chipselect;              // mm_interconnect_0:SECONDS_s1_chipselect -> SECONDS:chipselect
	wire  [31:0] mm_interconnect_0_seconds_s1_readdata;                // SECONDS:readdata -> mm_interconnect_0:SECONDS_s1_readdata
	wire   [1:0] mm_interconnect_0_seconds_s1_address;                 // mm_interconnect_0:SECONDS_s1_address -> SECONDS:address
	wire         mm_interconnect_0_seconds_s1_write;                   // mm_interconnect_0:SECONDS_s1_write -> SECONDS:write_n
	wire  [31:0] mm_interconnect_0_seconds_s1_writedata;               // mm_interconnect_0:SECONDS_s1_writedata -> SECONDS:writedata
	wire         mm_interconnect_0_minutes_s1_chipselect;              // mm_interconnect_0:MINUTES_s1_chipselect -> MINUTES:chipselect
	wire  [31:0] mm_interconnect_0_minutes_s1_readdata;                // MINUTES:readdata -> mm_interconnect_0:MINUTES_s1_readdata
	wire   [1:0] mm_interconnect_0_minutes_s1_address;                 // mm_interconnect_0:MINUTES_s1_address -> MINUTES:address
	wire         mm_interconnect_0_minutes_s1_write;                   // mm_interconnect_0:MINUTES_s1_write -> MINUTES:write_n
	wire  [31:0] mm_interconnect_0_minutes_s1_writedata;               // mm_interconnect_0:MINUTES_s1_writedata -> MINUTES:writedata
	wire         mm_interconnect_0_hours_s1_chipselect;                // mm_interconnect_0:HOURS_s1_chipselect -> HOURS:chipselect
	wire  [31:0] mm_interconnect_0_hours_s1_readdata;                  // HOURS:readdata -> mm_interconnect_0:HOURS_s1_readdata
	wire   [1:0] mm_interconnect_0_hours_s1_address;                   // mm_interconnect_0:HOURS_s1_address -> HOURS:address
	wire         mm_interconnect_0_hours_s1_write;                     // mm_interconnect_0:HOURS_s1_write -> HOURS:write_n
	wire  [31:0] mm_interconnect_0_hours_s1_writedata;                 // mm_interconnect_0:HOURS_s1_writedata -> HOURS:writedata
	wire         mm_interconnect_0_timercore_s1_chipselect;            // mm_interconnect_0:TimerCore_s1_chipselect -> TimerCore:chipselect
	wire  [15:0] mm_interconnect_0_timercore_s1_readdata;              // TimerCore:readdata -> mm_interconnect_0:TimerCore_s1_readdata
	wire   [2:0] mm_interconnect_0_timercore_s1_address;               // mm_interconnect_0:TimerCore_s1_address -> TimerCore:address
	wire         mm_interconnect_0_timercore_s1_write;                 // mm_interconnect_0:TimerCore_s1_write -> TimerCore:write_n
	wire  [15:0] mm_interconnect_0_timercore_s1_writedata;             // mm_interconnect_0:TimerCore_s1_writedata -> TimerCore:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;               // SWITCHES:readdata -> mm_interconnect_0:SWITCHES_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                // mm_interconnect_0:SWITCHES_s1_address -> SWITCHES:address
	wire         mm_interconnect_0_alarm_s1_chipselect;                // mm_interconnect_0:alarm_s1_chipselect -> alarm:chipselect
	wire  [31:0] mm_interconnect_0_alarm_s1_readdata;                  // alarm:readdata -> mm_interconnect_0:alarm_s1_readdata
	wire   [1:0] mm_interconnect_0_alarm_s1_address;                   // mm_interconnect_0:alarm_s1_address -> alarm:address
	wire         mm_interconnect_0_alarm_s1_write;                     // mm_interconnect_0:alarm_s1_write -> alarm:write_n
	wire  [31:0] mm_interconnect_0_alarm_s1_writedata;                 // mm_interconnect_0:alarm_s1_writedata -> alarm:writedata
	wire         irq_mapper_receiver0_irq;                             // UART:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // JTAG:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // TimerCore:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [BUTTONS:reset_n, CPU:reset_n, HOURS:reset_n, JTAG:rst_n, LEDs:reset_n, MINUTES:reset_n, RAM:reset, ROM:reset, SECONDS:reset_n, SWITCHES:reset_n, SysID:reset_n, TimerCore:reset_n, UART:reset, alarm:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                        // CPU:debug_reset_request -> rst_controller:reset_in1

	alarm_BUTTONS buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_export)                         // external_connection.export
	);

	alarm_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	alarm_HOURS hours (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_hours_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hours_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hours_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hours_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hours_s1_readdata),   //                    .readdata
		.out_port   (hours_export)                           // external_connection.export
	);

	alarm_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	alarm_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	alarm_HOURS minutes (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_minutes_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_minutes_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_minutes_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_minutes_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_minutes_s1_readdata),   //                    .readdata
		.out_port   (minutes_export)                           // external_connection.export
	);

	alarm_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	alarm_ROM rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	alarm_HOURS seconds (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_seconds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seconds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seconds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seconds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seconds_s1_readdata),   //                    .readdata
		.out_port   (seconds_export)                           // external_connection.export
	);

	alarm_SWITCHES switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	alarm_SysID sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	alarm_TimerCore timercore (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timercore_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timercore_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timercore_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timercore_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timercore_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                   //   irq.irq
	);

	alarm_UART uart (
		.clk        (clk_clk),                                              //                clk.clk
		.reset      (rst_controller_reset_out_reset),                       //              reset.reset
		.address    (mm_interconnect_0_uart_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_uart_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_uart_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_uart_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_uart_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_uart_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_uart_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver0_irq),                             //          interrupt.irq
		.UART_RXD   (uart_RXD),                                             // external_interface.export
		.UART_TXD   (uart_TXD)                                              //                   .export
	);

	alarm_alarm alarm (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_alarm_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_alarm_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_alarm_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_alarm_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_alarm_s1_readdata),   //                    .readdata
		.out_port   (alarm_export)                           // external_connection.export
	);

	alarm_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                           (clk_clk),                                              //                         CLK_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                              //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                          //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                           //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                                 //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                             //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                                //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                            //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                          //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                       //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                   //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                          //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                      //                                .readdata
		.alarm_s1_address                      (mm_interconnect_0_alarm_s1_address),                   //                        alarm_s1.address
		.alarm_s1_write                        (mm_interconnect_0_alarm_s1_write),                     //                                .write
		.alarm_s1_readdata                     (mm_interconnect_0_alarm_s1_readdata),                  //                                .readdata
		.alarm_s1_writedata                    (mm_interconnect_0_alarm_s1_writedata),                 //                                .writedata
		.alarm_s1_chipselect                   (mm_interconnect_0_alarm_s1_chipselect),                //                                .chipselect
		.BUTTONS_s1_address                    (mm_interconnect_0_buttons_s1_address),                 //                      BUTTONS_s1.address
		.BUTTONS_s1_readdata                   (mm_interconnect_0_buttons_s1_readdata),                //                                .readdata
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),        //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                .debugaccess
		.HOURS_s1_address                      (mm_interconnect_0_hours_s1_address),                   //                        HOURS_s1.address
		.HOURS_s1_write                        (mm_interconnect_0_hours_s1_write),                     //                                .write
		.HOURS_s1_readdata                     (mm_interconnect_0_hours_s1_readdata),                  //                                .readdata
		.HOURS_s1_writedata                    (mm_interconnect_0_hours_s1_writedata),                 //                                .writedata
		.HOURS_s1_chipselect                   (mm_interconnect_0_hours_s1_chipselect),                //                                .chipselect
		.JTAG_avalon_jtag_slave_address        (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //          JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write          (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                .write
		.JTAG_avalon_jtag_slave_read           (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                .read
		.JTAG_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                .readdata
		.JTAG_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                .writedata
		.JTAG_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.JTAG_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                .chipselect
		.LEDs_s1_address                       (mm_interconnect_0_leds_s1_address),                    //                         LEDs_s1.address
		.LEDs_s1_write                         (mm_interconnect_0_leds_s1_write),                      //                                .write
		.LEDs_s1_readdata                      (mm_interconnect_0_leds_s1_readdata),                   //                                .readdata
		.LEDs_s1_writedata                     (mm_interconnect_0_leds_s1_writedata),                  //                                .writedata
		.LEDs_s1_chipselect                    (mm_interconnect_0_leds_s1_chipselect),                 //                                .chipselect
		.MINUTES_s1_address                    (mm_interconnect_0_minutes_s1_address),                 //                      MINUTES_s1.address
		.MINUTES_s1_write                      (mm_interconnect_0_minutes_s1_write),                   //                                .write
		.MINUTES_s1_readdata                   (mm_interconnect_0_minutes_s1_readdata),                //                                .readdata
		.MINUTES_s1_writedata                  (mm_interconnect_0_minutes_s1_writedata),               //                                .writedata
		.MINUTES_s1_chipselect                 (mm_interconnect_0_minutes_s1_chipselect),              //                                .chipselect
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                     //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                       //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                    //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                   //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),                  //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),                  //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                       //                                .clken
		.ROM_s1_address                        (mm_interconnect_0_rom_s1_address),                     //                          ROM_s1.address
		.ROM_s1_write                          (mm_interconnect_0_rom_s1_write),                       //                                .write
		.ROM_s1_readdata                       (mm_interconnect_0_rom_s1_readdata),                    //                                .readdata
		.ROM_s1_writedata                      (mm_interconnect_0_rom_s1_writedata),                   //                                .writedata
		.ROM_s1_byteenable                     (mm_interconnect_0_rom_s1_byteenable),                  //                                .byteenable
		.ROM_s1_chipselect                     (mm_interconnect_0_rom_s1_chipselect),                  //                                .chipselect
		.ROM_s1_clken                          (mm_interconnect_0_rom_s1_clken),                       //                                .clken
		.ROM_s1_debugaccess                    (mm_interconnect_0_rom_s1_debugaccess),                 //                                .debugaccess
		.SECONDS_s1_address                    (mm_interconnect_0_seconds_s1_address),                 //                      SECONDS_s1.address
		.SECONDS_s1_write                      (mm_interconnect_0_seconds_s1_write),                   //                                .write
		.SECONDS_s1_readdata                   (mm_interconnect_0_seconds_s1_readdata),                //                                .readdata
		.SECONDS_s1_writedata                  (mm_interconnect_0_seconds_s1_writedata),               //                                .writedata
		.SECONDS_s1_chipselect                 (mm_interconnect_0_seconds_s1_chipselect),              //                                .chipselect
		.SWITCHES_s1_address                   (mm_interconnect_0_switches_s1_address),                //                     SWITCHES_s1.address
		.SWITCHES_s1_readdata                  (mm_interconnect_0_switches_s1_readdata),               //                                .readdata
		.SysID_control_slave_address           (mm_interconnect_0_sysid_control_slave_address),        //             SysID_control_slave.address
		.SysID_control_slave_readdata          (mm_interconnect_0_sysid_control_slave_readdata),       //                                .readdata
		.TimerCore_s1_address                  (mm_interconnect_0_timercore_s1_address),               //                    TimerCore_s1.address
		.TimerCore_s1_write                    (mm_interconnect_0_timercore_s1_write),                 //                                .write
		.TimerCore_s1_readdata                 (mm_interconnect_0_timercore_s1_readdata),              //                                .readdata
		.TimerCore_s1_writedata                (mm_interconnect_0_timercore_s1_writedata),             //                                .writedata
		.TimerCore_s1_chipselect               (mm_interconnect_0_timercore_s1_chipselect),            //                                .chipselect
		.UART_avalon_rs232_slave_address       (mm_interconnect_0_uart_avalon_rs232_slave_address),    //         UART_avalon_rs232_slave.address
		.UART_avalon_rs232_slave_write         (mm_interconnect_0_uart_avalon_rs232_slave_write),      //                                .write
		.UART_avalon_rs232_slave_read          (mm_interconnect_0_uart_avalon_rs232_slave_read),       //                                .read
		.UART_avalon_rs232_slave_readdata      (mm_interconnect_0_uart_avalon_rs232_slave_readdata),   //                                .readdata
		.UART_avalon_rs232_slave_writedata     (mm_interconnect_0_uart_avalon_rs232_slave_writedata),  //                                .writedata
		.UART_avalon_rs232_slave_byteenable    (mm_interconnect_0_uart_avalon_rs232_slave_byteenable), //                                .byteenable
		.UART_avalon_rs232_slave_chipselect    (mm_interconnect_0_uart_avalon_rs232_slave_chipselect)  //                                .chipselect
	);

	alarm_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
