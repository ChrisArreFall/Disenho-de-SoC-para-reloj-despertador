// NIOS_SoC.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NIOS_SoC (
		input  wire [3:0] btn_export,    //    btn.export
		input  wire       clk_clk,       //    clk.clk
		output wire [6:0] hex0_export,   //   hex0.export
		output wire [6:0] hex1_export,   //   hex1.export
		output wire [6:0] hex2_export,   //   hex2.export
		output wire [6:0] hex3_export,   //   hex3.export
		output wire [6:0] hex4_export,   //   hex4.export
		output wire [6:0] hex5_export,   //   hex5.export
		input  wire       reset_reset_n, //  reset.reset_n
		output wire       timer_export,  //  timer.export
		input  wire       uartpc_rxd,    // uartpc.rxd
		output wire       uartpc_txd     //       .txd
	);

	wire  [31:0] nios_data_master_readdata;                          // mm_interconnect_0:NIOS_data_master_readdata -> NIOS:d_readdata
	wire         nios_data_master_waitrequest;                       // mm_interconnect_0:NIOS_data_master_waitrequest -> NIOS:d_waitrequest
	wire         nios_data_master_debugaccess;                       // NIOS:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_data_master_debugaccess
	wire  [13:0] nios_data_master_address;                           // NIOS:d_address -> mm_interconnect_0:NIOS_data_master_address
	wire   [3:0] nios_data_master_byteenable;                        // NIOS:d_byteenable -> mm_interconnect_0:NIOS_data_master_byteenable
	wire         nios_data_master_read;                              // NIOS:d_read -> mm_interconnect_0:NIOS_data_master_read
	wire         nios_data_master_write;                             // NIOS:d_write -> mm_interconnect_0:NIOS_data_master_write
	wire  [31:0] nios_data_master_writedata;                         // NIOS:d_writedata -> mm_interconnect_0:NIOS_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                   // mm_interconnect_0:NIOS_instruction_master_readdata -> NIOS:i_readdata
	wire         nios_instruction_master_waitrequest;                // mm_interconnect_0:NIOS_instruction_master_waitrequest -> NIOS:i_waitrequest
	wire  [13:0] nios_instruction_master_address;                    // NIOS:i_address -> mm_interconnect_0:NIOS_instruction_master_address
	wire         nios_instruction_master_read;                       // NIOS:i_read -> mm_interconnect_0:NIOS_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;    // NIOS:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest; // NIOS:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess; // mm_interconnect_0:NIOS_debug_mem_slave_debugaccess -> NIOS:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;     // mm_interconnect_0:NIOS_debug_mem_slave_address -> NIOS:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;        // mm_interconnect_0:NIOS_debug_mem_slave_read -> NIOS:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;  // mm_interconnect_0:NIOS_debug_mem_slave_byteenable -> NIOS:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;       // mm_interconnect_0:NIOS_debug_mem_slave_write -> NIOS:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;   // mm_interconnect_0:NIOS_debug_mem_slave_writedata -> NIOS:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;             // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;               // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [9:0] mm_interconnect_0_memory_s1_address;                // mm_interconnect_0:memory_s1_address -> memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;             // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                  // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;              // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                  // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_segment0_s1_chipselect;           // mm_interconnect_0:Segment0_s1_chipselect -> Segment0:chipselect
	wire  [31:0] mm_interconnect_0_segment0_s1_readdata;             // Segment0:readdata -> mm_interconnect_0:Segment0_s1_readdata
	wire   [1:0] mm_interconnect_0_segment0_s1_address;              // mm_interconnect_0:Segment0_s1_address -> Segment0:address
	wire         mm_interconnect_0_segment0_s1_write;                // mm_interconnect_0:Segment0_s1_write -> Segment0:write_n
	wire  [31:0] mm_interconnect_0_segment0_s1_writedata;            // mm_interconnect_0:Segment0_s1_writedata -> Segment0:writedata
	wire  [31:0] mm_interconnect_0_button_s1_readdata;               // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_segment1_s1_chipselect;           // mm_interconnect_0:Segment1_s1_chipselect -> Segment1:chipselect
	wire  [31:0] mm_interconnect_0_segment1_s1_readdata;             // Segment1:readdata -> mm_interconnect_0:Segment1_s1_readdata
	wire   [1:0] mm_interconnect_0_segment1_s1_address;              // mm_interconnect_0:Segment1_s1_address -> Segment1:address
	wire         mm_interconnect_0_segment1_s1_write;                // mm_interconnect_0:Segment1_s1_write -> Segment1:write_n
	wire  [31:0] mm_interconnect_0_segment1_s1_writedata;            // mm_interconnect_0:Segment1_s1_writedata -> Segment1:writedata
	wire         mm_interconnect_0_segment3_s1_chipselect;           // mm_interconnect_0:Segment3_s1_chipselect -> Segment3:chipselect
	wire  [31:0] mm_interconnect_0_segment3_s1_readdata;             // Segment3:readdata -> mm_interconnect_0:Segment3_s1_readdata
	wire   [1:0] mm_interconnect_0_segment3_s1_address;              // mm_interconnect_0:Segment3_s1_address -> Segment3:address
	wire         mm_interconnect_0_segment3_s1_write;                // mm_interconnect_0:Segment3_s1_write -> Segment3:write_n
	wire  [31:0] mm_interconnect_0_segment3_s1_writedata;            // mm_interconnect_0:Segment3_s1_writedata -> Segment3:writedata
	wire         mm_interconnect_0_segment2_s1_chipselect;           // mm_interconnect_0:Segment2_s1_chipselect -> Segment2:chipselect
	wire  [31:0] mm_interconnect_0_segment2_s1_readdata;             // Segment2:readdata -> mm_interconnect_0:Segment2_s1_readdata
	wire   [1:0] mm_interconnect_0_segment2_s1_address;              // mm_interconnect_0:Segment2_s1_address -> Segment2:address
	wire         mm_interconnect_0_segment2_s1_write;                // mm_interconnect_0:Segment2_s1_write -> Segment2:write_n
	wire  [31:0] mm_interconnect_0_segment2_s1_writedata;            // mm_interconnect_0:Segment2_s1_writedata -> Segment2:writedata
	wire         mm_interconnect_0_segment4_s1_chipselect;           // mm_interconnect_0:Segment4_s1_chipselect -> Segment4:chipselect
	wire  [31:0] mm_interconnect_0_segment4_s1_readdata;             // Segment4:readdata -> mm_interconnect_0:Segment4_s1_readdata
	wire   [1:0] mm_interconnect_0_segment4_s1_address;              // mm_interconnect_0:Segment4_s1_address -> Segment4:address
	wire         mm_interconnect_0_segment4_s1_write;                // mm_interconnect_0:Segment4_s1_write -> Segment4:write_n
	wire  [31:0] mm_interconnect_0_segment4_s1_writedata;            // mm_interconnect_0:Segment4_s1_writedata -> Segment4:writedata
	wire         mm_interconnect_0_segment5_s1_chipselect;           // mm_interconnect_0:Segment5_s1_chipselect -> Segment5:chipselect
	wire  [31:0] mm_interconnect_0_segment5_s1_readdata;             // Segment5:readdata -> mm_interconnect_0:Segment5_s1_readdata
	wire   [1:0] mm_interconnect_0_segment5_s1_address;              // mm_interconnect_0:Segment5_s1_address -> Segment5:address
	wire         mm_interconnect_0_segment5_s1_write;                // mm_interconnect_0:Segment5_s1_write -> Segment5:write_n
	wire  [31:0] mm_interconnect_0_segment5_s1_writedata;            // mm_interconnect_0:Segment5_s1_writedata -> Segment5:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;              // mm_interconnect_0:Timer_s1_chipselect -> Timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                // Timer:readdata -> mm_interconnect_0:Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                 // mm_interconnect_0:Timer_s1_address -> Timer:address
	wire         mm_interconnect_0_timer_s1_write;                   // mm_interconnect_0:Timer_s1_write -> Timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;               // mm_interconnect_0:Timer_s1_writedata -> Timer:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;               // mm_interconnect_0:UART_s1_chipselect -> UART:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                 // UART:readdata -> mm_interconnect_0:UART_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                  // mm_interconnect_0:UART_s1_address -> UART:address
	wire         mm_interconnect_0_uart_s1_read;                     // mm_interconnect_0:UART_s1_read -> UART:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;            // mm_interconnect_0:UART_s1_begintransfer -> UART:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                    // mm_interconnect_0:UART_s1_write -> UART:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                // mm_interconnect_0:UART_s1_writedata -> UART:writedata
	wire         irq_mapper_receiver0_irq;                           // Timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                           // UART:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_irq_irq;                                       // irq_mapper:sender_irq -> NIOS:irq
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [NIOS:reset_n, Segment0:reset_n, Segment1:reset_n, Segment2:reset_n, Segment3:reset_n, Segment4:reset_n, Segment5:reset_n, Timer:reset_n, UART:reset_n, irq_mapper:reset, memory:reset, mm_interconnect_0:NIOS_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [NIOS:reset_req, memory:reset_req, rst_translator:reset_req_in]
	wire         nios_debug_reset_request_reset;                     // NIOS:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> [button:reset_n, mm_interconnect_0:button_reset_reset_bridge_in_reset_reset]

	NIOS_SoC_NIOS nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	NIOS_SoC_Segment0 segment0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment0_s1_readdata),   //                    .readdata
		.out_port   (hex0_export)                               // external_connection.export
	);

	NIOS_SoC_Segment0 segment1 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment1_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                               // external_connection.export
	);

	NIOS_SoC_Segment0 segment2 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment2_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                               // external_connection.export
	);

	NIOS_SoC_Segment0 segment3 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment3_s1_readdata),   //                    .readdata
		.out_port   (hex3_export)                               // external_connection.export
	);

	NIOS_SoC_Segment0 segment4 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment4_s1_readdata),   //                    .readdata
		.out_port   (hex4_export)                               // external_connection.export
	);

	NIOS_SoC_Segment0 segment5 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_segment5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segment5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segment5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segment5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segment5_s1_readdata),   //                    .readdata
		.out_port   (hex5_export)                               // external_connection.export
	);

	NIOS_SoC_Timer timer (
		.clk           (clk_clk),                               //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),       //         reset.reset_n
		.address       (mm_interconnect_0_timer_s1_address),    //            s1.address
		.writedata     (mm_interconnect_0_timer_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_0_timer_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_0_timer_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_0_timer_s1_write),     //              .write_n
		.irq           (irq_mapper_receiver0_irq),              //           irq.irq
		.timeout_pulse (timer_export)                           // external_port.export
	);

	NIOS_SoC_UART uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uartpc_rxd),                              // external_connection.export
		.txd           (uartpc_txd),                              //                    .export
		.irq           (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	NIOS_SoC_button button (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_s1_readdata), //                    .readdata
		.in_port  (btn_export)                            // external_connection.export
	);

	NIOS_SoC_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	NIOS_SoC_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (clk_clk),                                            //                            clk_clk.clk
		.button_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                 // button_reset_reset_bridge_in_reset.reset
		.NIOS_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                     //   NIOS_reset_reset_bridge_in_reset.reset
		.NIOS_data_master_address                 (nios_data_master_address),                           //                   NIOS_data_master.address
		.NIOS_data_master_waitrequest             (nios_data_master_waitrequest),                       //                                   .waitrequest
		.NIOS_data_master_byteenable              (nios_data_master_byteenable),                        //                                   .byteenable
		.NIOS_data_master_read                    (nios_data_master_read),                              //                                   .read
		.NIOS_data_master_readdata                (nios_data_master_readdata),                          //                                   .readdata
		.NIOS_data_master_write                   (nios_data_master_write),                             //                                   .write
		.NIOS_data_master_writedata               (nios_data_master_writedata),                         //                                   .writedata
		.NIOS_data_master_debugaccess             (nios_data_master_debugaccess),                       //                                   .debugaccess
		.NIOS_instruction_master_address          (nios_instruction_master_address),                    //            NIOS_instruction_master.address
		.NIOS_instruction_master_waitrequest      (nios_instruction_master_waitrequest),                //                                   .waitrequest
		.NIOS_instruction_master_read             (nios_instruction_master_read),                       //                                   .read
		.NIOS_instruction_master_readdata         (nios_instruction_master_readdata),                   //                                   .readdata
		.button_s1_address                        (mm_interconnect_0_button_s1_address),                //                          button_s1.address
		.button_s1_readdata                       (mm_interconnect_0_button_s1_readdata),               //                                   .readdata
		.memory_s1_address                        (mm_interconnect_0_memory_s1_address),                //                          memory_s1.address
		.memory_s1_write                          (mm_interconnect_0_memory_s1_write),                  //                                   .write
		.memory_s1_readdata                       (mm_interconnect_0_memory_s1_readdata),               //                                   .readdata
		.memory_s1_writedata                      (mm_interconnect_0_memory_s1_writedata),              //                                   .writedata
		.memory_s1_byteenable                     (mm_interconnect_0_memory_s1_byteenable),             //                                   .byteenable
		.memory_s1_chipselect                     (mm_interconnect_0_memory_s1_chipselect),             //                                   .chipselect
		.memory_s1_clken                          (mm_interconnect_0_memory_s1_clken),                  //                                   .clken
		.NIOS_debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //               NIOS_debug_mem_slave.address
		.NIOS_debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                                   .write
		.NIOS_debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                                   .read
		.NIOS_debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                                   .readdata
		.NIOS_debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                                   .writedata
		.NIOS_debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                                   .byteenable
		.NIOS_debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                                   .waitrequest
		.NIOS_debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                                   .debugaccess
		.Segment0_s1_address                      (mm_interconnect_0_segment0_s1_address),              //                        Segment0_s1.address
		.Segment0_s1_write                        (mm_interconnect_0_segment0_s1_write),                //                                   .write
		.Segment0_s1_readdata                     (mm_interconnect_0_segment0_s1_readdata),             //                                   .readdata
		.Segment0_s1_writedata                    (mm_interconnect_0_segment0_s1_writedata),            //                                   .writedata
		.Segment0_s1_chipselect                   (mm_interconnect_0_segment0_s1_chipselect),           //                                   .chipselect
		.Segment1_s1_address                      (mm_interconnect_0_segment1_s1_address),              //                        Segment1_s1.address
		.Segment1_s1_write                        (mm_interconnect_0_segment1_s1_write),                //                                   .write
		.Segment1_s1_readdata                     (mm_interconnect_0_segment1_s1_readdata),             //                                   .readdata
		.Segment1_s1_writedata                    (mm_interconnect_0_segment1_s1_writedata),            //                                   .writedata
		.Segment1_s1_chipselect                   (mm_interconnect_0_segment1_s1_chipselect),           //                                   .chipselect
		.Segment2_s1_address                      (mm_interconnect_0_segment2_s1_address),              //                        Segment2_s1.address
		.Segment2_s1_write                        (mm_interconnect_0_segment2_s1_write),                //                                   .write
		.Segment2_s1_readdata                     (mm_interconnect_0_segment2_s1_readdata),             //                                   .readdata
		.Segment2_s1_writedata                    (mm_interconnect_0_segment2_s1_writedata),            //                                   .writedata
		.Segment2_s1_chipselect                   (mm_interconnect_0_segment2_s1_chipselect),           //                                   .chipselect
		.Segment3_s1_address                      (mm_interconnect_0_segment3_s1_address),              //                        Segment3_s1.address
		.Segment3_s1_write                        (mm_interconnect_0_segment3_s1_write),                //                                   .write
		.Segment3_s1_readdata                     (mm_interconnect_0_segment3_s1_readdata),             //                                   .readdata
		.Segment3_s1_writedata                    (mm_interconnect_0_segment3_s1_writedata),            //                                   .writedata
		.Segment3_s1_chipselect                   (mm_interconnect_0_segment3_s1_chipselect),           //                                   .chipselect
		.Segment4_s1_address                      (mm_interconnect_0_segment4_s1_address),              //                        Segment4_s1.address
		.Segment4_s1_write                        (mm_interconnect_0_segment4_s1_write),                //                                   .write
		.Segment4_s1_readdata                     (mm_interconnect_0_segment4_s1_readdata),             //                                   .readdata
		.Segment4_s1_writedata                    (mm_interconnect_0_segment4_s1_writedata),            //                                   .writedata
		.Segment4_s1_chipselect                   (mm_interconnect_0_segment4_s1_chipselect),           //                                   .chipselect
		.Segment5_s1_address                      (mm_interconnect_0_segment5_s1_address),              //                        Segment5_s1.address
		.Segment5_s1_write                        (mm_interconnect_0_segment5_s1_write),                //                                   .write
		.Segment5_s1_readdata                     (mm_interconnect_0_segment5_s1_readdata),             //                                   .readdata
		.Segment5_s1_writedata                    (mm_interconnect_0_segment5_s1_writedata),            //                                   .writedata
		.Segment5_s1_chipselect                   (mm_interconnect_0_segment5_s1_chipselect),           //                                   .chipselect
		.Timer_s1_address                         (mm_interconnect_0_timer_s1_address),                 //                           Timer_s1.address
		.Timer_s1_write                           (mm_interconnect_0_timer_s1_write),                   //                                   .write
		.Timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),                //                                   .readdata
		.Timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),               //                                   .writedata
		.Timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect),              //                                   .chipselect
		.UART_s1_address                          (mm_interconnect_0_uart_s1_address),                  //                            UART_s1.address
		.UART_s1_write                            (mm_interconnect_0_uart_s1_write),                    //                                   .write
		.UART_s1_read                             (mm_interconnect_0_uart_s1_read),                     //                                   .read
		.UART_s1_readdata                         (mm_interconnect_0_uart_s1_readdata),                 //                                   .readdata
		.UART_s1_writedata                        (mm_interconnect_0_uart_s1_writedata),                //                                   .writedata
		.UART_s1_begintransfer                    (mm_interconnect_0_uart_s1_begintransfer),            //                                   .begintransfer
		.UART_s1_chipselect                       (mm_interconnect_0_uart_s1_chipselect)                //                                   .chipselect
	);

	NIOS_SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_debug_reset_request_reset),     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
